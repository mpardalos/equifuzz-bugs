module spec(out);
  output wire  [40:0] out;
  assign out = 41'b000000000000000000000000000000000000000000;
endmodule
