module spec(out);
  output wire signed [42:0] out;
  assign out = 43'b0000000000000000000000000000000000000000000;
endmodule
