module spec(out);
  output wire  [40:0] out;
  assign out = 41'b00000000000000000000000000000000000000000;
endmodule
