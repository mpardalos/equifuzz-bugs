module spec (out);
  output wire signed [15:0] out;
  assign out = 16'b0000000100000000;
endmodule
