module spec (out);
  output wire signed [7:0] out;
  assign out = 8'b0000000100000000;
endmodule
